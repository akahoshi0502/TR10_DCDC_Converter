* Extracted by KLayout

.SUBCKT SA_VCO_TOP VDD BIAS_IN OUT VSS
X$1 VDD \$4 BIAS_IN VSS SA_VCO
X$2 VDD \$4 OUT VSS SA_DFF_Counter_8
.ENDS SA_VCO_TOP

.SUBCKT SA_VCO VDD OUT \$8 VSS
X$1 VDD \$I287 \$2 \$9 VSS SA_VCO_INV
X$2 VDD \$2 \$I269 \$9 VSS SA_VCO_INV
X$16 VDD \$I255 \$I287 \$9 VSS SA_VCO_INV
X$25 VDD \$I256 \$I255 \$9 VSS SA_VCO_INV
X$34 VDD \$I257 \$I256 \$9 VSS SA_VCO_INV
X$43 VDD \$I258 \$I257 \$9 VSS SA_VCO_INV
X$52 VDD \$I259 \$I258 \$9 VSS SA_VCO_INV
X$61 VDD \$I260 \$I259 \$9 VSS SA_VCO_INV
X$70 VDD \$I261 \$I260 \$9 VSS SA_VCO_INV
X$79 VDD OUT \$I261 \$9 VSS SA_VCO_INV
X$92 VDD \$I263 OUT \$9 VSS SA_VCO_INV
X$101 VDD \$I264 \$I263 \$9 VSS SA_VCO_INV
X$110 VDD \$I265 \$I264 \$9 VSS SA_VCO_INV
X$119 VDD \$I266 \$I265 \$9 VSS SA_VCO_INV
X$128 VDD \$I267 \$I266 \$9 VSS SA_VCO_INV
X$137 VDD \$I268 \$I267 \$9 VSS SA_VCO_INV
X$146 VDD \$I269 \$I268 \$9 VSS SA_VCO_INV
M$1 VSS VSS VSS VSS NCHOR1EX L=1U W=20U AS=38P AD=38P PS=60U PD=60U
M$2 \$9 \$8 VSS VSS NCHOR1EX L=1U W=8U AS=8P AD=8P PS=16U PD=16U
M$7 VDD VDD VDD VDD PCHOR1EX L=1U W=16U AS=32P AD=32P PS=48U PD=48U
.ENDS SA_VCO

.SUBCKT SA_DFF_Counter_8 VDD IN OUT VSS
X$1 \$I15 \$I1 VDD VSS SA_DFF_Counter
X$2 IN \$I15 VDD VSS SA_DFF_Counter
X$3 \$I1 \$I2 VDD VSS SA_DFF_Counter
X$4 \$I2 \$I3 VDD VSS SA_DFF_Counter
X$5 \$I3 \$I4 VDD VSS SA_DFF_Counter
X$6 \$I4 \$I5 VDD VSS SA_DFF_Counter
X$7 \$I5 \$I6 VDD VSS SA_DFF_Counter
X$8 \$I6 OUT VDD VSS SA_DFF_Counter
.ENDS SA_DFF_Counter_8

.SUBCKT SA_VCO_INV VDD OUT IN nchSource VSS
M$1 VSS OUT VSS VSS NCHOR1EX L=3U W=6U AS=12P AD=12P PS=16U PD=16U
M$2 OUT IN VDD VDD PCHOR1EX L=1U W=16U AS=20P AD=20P PS=30U PD=30U
M$6 OUT IN nchSource VSS NCHOR1EX L=1U W=8U AS=12P AD=12P PS=18U PD=18U
.ENDS SA_VCO_INV

.SUBCKT SA_DFF_Counter IN OUT VDD VSS
X$1 IN \$5 \$5 OUT VDD VSS dff1
.ENDS SA_DFF_Counter

.SUBCKT dff1 CK D QB Q VDD VSS
M$1 VDD \$11 QB VDD PCHOR1EX L=1U W=6U AS=12P AD=6P PS=16U PD=8U
M$2 Q QB VDD VDD PCHOR1EX L=1U W=6U AS=6P AD=12P PS=8U PD=16U
M$3 \$69 \$8 VDD VDD PCHOR1EX L=1U W=6U AS=12P AD=3P PS=16U PD=7U
M$4 \$38 \$4 \$69 VDD PCHOR1EX L=1U W=6U AS=3P AD=6P PS=7U PD=8U
M$5 \$70 \$2 \$38 VDD PCHOR1EX L=1U W=6U AS=6P AD=3P PS=8U PD=7U
M$6 VDD \$11 \$70 VDD PCHOR1EX L=1U W=6U AS=3P AD=6P PS=7U PD=8U
M$7 \$11 \$38 VDD VDD PCHOR1EX L=1U W=6U AS=6P AD=12P PS=8U PD=16U
M$8 VDD CK \$2 VDD PCHOR1EX L=1U W=6U AS=12P AD=6P PS=16U PD=8U
M$9 \$4 \$2 VDD VDD PCHOR1EX L=1U W=6U AS=6P AD=12P PS=8U PD=16U
M$10 \$63 D VDD VDD PCHOR1EX L=1U W=6U AS=12P AD=3P PS=16U PD=7U
M$11 \$7 \$2 \$63 VDD PCHOR1EX L=1U W=6U AS=3P AD=6P PS=7U PD=8U
M$12 \$65 \$4 \$7 VDD PCHOR1EX L=1U W=6U AS=6P AD=3P PS=8U PD=7U
M$13 VDD \$8 \$65 VDD PCHOR1EX L=1U W=6U AS=3P AD=6P PS=7U PD=8U
M$14 \$8 \$7 VDD VDD PCHOR1EX L=1U W=6U AS=6P AD=12P PS=8U PD=16U
M$15 VSS \$11 QB VSS NCHOR1EX L=1U W=2U AS=4P AD=2P PS=8U PD=4U
M$16 Q QB VSS VSS NCHOR1EX L=1U W=2U AS=2P AD=4P PS=4U PD=8U
M$17 \$36 \$8 VSS VSS NCHOR1EX L=1U W=2U AS=4P AD=1P PS=8U PD=3U
M$18 \$38 \$2 \$36 VSS NCHOR1EX L=1U W=2U AS=1P AD=2P PS=3U PD=4U
M$19 \$41 \$4 \$38 VSS NCHOR1EX L=1U W=2U AS=2P AD=1P PS=4U PD=3U
M$20 VSS \$11 \$41 VSS NCHOR1EX L=1U W=2U AS=1P AD=2P PS=3U PD=4U
M$21 \$11 \$38 VSS VSS NCHOR1EX L=1U W=2U AS=2P AD=4P PS=4U PD=8U
M$22 VSS CK \$2 VSS NCHOR1EX L=1U W=2U AS=4P AD=2P PS=8U PD=4U
M$23 \$4 \$2 VSS VSS NCHOR1EX L=1U W=2U AS=2P AD=4P PS=4U PD=8U
M$24 \$22 D VSS VSS NCHOR1EX L=1U W=2U AS=4P AD=1P PS=8U PD=3U
M$25 \$7 \$4 \$22 VSS NCHOR1EX L=1U W=2U AS=1P AD=2P PS=3U PD=4U
M$26 \$26 \$2 \$7 VSS NCHOR1EX L=1U W=2U AS=2P AD=1P PS=4U PD=3U
M$27 VSS \$8 \$26 VSS NCHOR1EX L=1U W=2U AS=1P AD=2P PS=3U PD=4U
M$28 \$8 \$7 VSS VSS NCHOR1EX L=1U W=2U AS=2P AD=4P PS=4U PD=8U
.ENDS dff1
