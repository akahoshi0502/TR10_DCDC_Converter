* Extracted by KLayout

.SUBCKT SA_VCO_DECAP_B VDD VSS
C$1 VSS VDD 7.9866e-13 POLY_CAP
.ENDS SA_VCO_DECAP_B
